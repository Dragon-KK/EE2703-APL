.circuit # An empty circuit
.end